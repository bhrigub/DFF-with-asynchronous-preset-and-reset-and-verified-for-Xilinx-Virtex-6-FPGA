library verilog;
use verilog.vl_types.all;
entity tbd is
end tbd;
